module hw1(
	input CLK_50M,
	input RESET_N,
	
);

	

endmodule 