module tx_time_gen(
	input CLK,
	input reset,
	output reg tick
);

		reg [] counter;
		
		always@(posedge CLK,negedge reset)begin
			
		end

endmodule