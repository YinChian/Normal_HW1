module hw1(
	input CLK_50M,
	input RESET_N,
	input [7:0] write_data,
	input write,
	output uart_txd,
	
	input uart_rxd,
	output read_error,
	output read_complete,
	output [7:0] read_value
);

	

endmodule 